module sec_ded_daec_decoder_64(
  input  logic        clk,
  input  logic[63:0]  data_i,
  input  logic[7:0]   ecc_i,
  output logic[63:0]  corrected_data_o,
  output logic        uncorrectable_error_o
);

  logic[7:0]  syndrome;
  logic[7:0]  syndrome_next;
  logic[63:0] data_next;
  logic[63:0] error_mask;

  //  row0: 0 3 5 7 8 9 11 13 14 17 19 22 25 30 32 33 37 40 41 44 48 49 51 56 57 58
  //  row1: 0 2 3 4 7 8 14 16 18 21 24 29 31 32 36 39 40 43 47 48 50 55 56 57 63
  //  row2: 1 2 4 6 8 10 11 12 14 16 17 20 23 28 30 31 35 38 39 42 46 47 49 54 55 56 62 63
  //  row3: 0 1 2 3 5 6 9 11 12 15 16 19 22 24 27 29 30 34 37 38 41 45 46 48 53 54 61 62 63
  //  row4: 0 3 5 6 10 11 12 13 15 16 18 21 23 26 28 29 33 36 37 40 44 45 52 53 55 60 61 62
  //  row5: 0 1 2 4 5 8 9 10 11 12 13 15 16 17 20 22 25 27 28 32 35 36 43 44 47 51 52 54 59 60 61
  //  row6: 1 2 4 6 7 9 10 12 13 14 15 19 21 24 26 27 34 35 39 42 43 46 50 51 53 58 59 60
  //  row7: 1 3 4 5 6 8 9 10 13 14 15 18 20 23 25 26 31 33 34 38 41 42 45 49 50 52 57 58 59

  assign syndrome[0] = ecc_i[0]^data_i[0]^data_i[3]^data_i[5]^data_i[7]^data_i[8]^data_i[9]^data_i[11]^data_i[13]^data_i[14]^data_i[17]^data_i[19]^data_i[22]^data_i[25]^data_i[30]^data_i[32]^data_i[33]^data_i[37]^data_i[40]^data_i[41]^data_i[44]^data_i[48]^data_i[49]^data_i[51]^data_i[56]^data_i[57]^data_i[58];
  assign syndrome[1] = ecc_i[1]^data_i[0]^data_i[2]^data_i[3]^data_i[4]^data_i[7]^data_i[8]^data_i[14]^data_i[16]^data_i[18]^data_i[21]^data_i[24]^data_i[29]^data_i[31]^data_i[32]^data_i[36]^data_i[39]^data_i[40]^data_i[43]^data_i[47]^data_i[48]^data_i[50]^data_i[55]^data_i[56]^data_i[57]^data_i[63];
  assign syndrome[2] = ecc_i[2]^data_i[1]^data_i[2]^data_i[4]^data_i[6]^data_i[8]^data_i[10]^data_i[11]^data_i[12]^data_i[14]^data_i[16]^data_i[17]^data_i[20]^data_i[23]^data_i[28]^data_i[30]^data_i[31]^data_i[35]^data_i[38]^data_i[39]^data_i[42]^data_i[46]^data_i[47]^data_i[49]^data_i[54]^data_i[55]^data_i[56]^data_i[62]^data_i[63];
  assign syndrome[3] = ecc_i[3]^data_i[0]^data_i[1]^data_i[2]^data_i[3]^data_i[5]^data_i[6]^data_i[9]^data_i[11]^data_i[12]^data_i[15]^data_i[16]^data_i[19]^data_i[22]^data_i[24]^data_i[27]^data_i[29]^data_i[30]^data_i[34]^data_i[37]^data_i[38]^data_i[41]^data_i[45]^data_i[46]^data_i[48]^data_i[53]^data_i[54]^data_i[61]^data_i[62]^data_i[63];
  assign syndrome[4] = ecc_i[4]^data_i[0]^data_i[3]^data_i[5]^data_i[6]^data_i[10]^data_i[11]^data_i[12]^data_i[13]^data_i[15]^data_i[16]^data_i[18]^data_i[21]^data_i[23]^data_i[26]^data_i[28]^data_i[29]^data_i[33]^data_i[36]^data_i[37]^data_i[40]^data_i[44]^data_i[45]^data_i[52]^data_i[53]^data_i[55]^data_i[60]^data_i[61]^data_i[62];
  assign syndrome[5] = ecc_i[5]^data_i[0]^data_i[1]^data_i[2]^data_i[4]^data_i[5]^data_i[8]^data_i[9]^data_i[10]^data_i[11]^data_i[12]^data_i[13]^data_i[15]^data_i[16]^data_i[17]^data_i[20]^data_i[22]^data_i[25]^data_i[27]^data_i[28]^data_i[32]^data_i[35]^data_i[36]^data_i[43]^data_i[44]^data_i[47]^data_i[51]^data_i[52]^data_i[54]^data_i[59]^data_i[60]^data_i[61];
  assign syndrome[6] = ecc_i[6]^data_i[1]^data_i[2]^data_i[4]^data_i[6]^data_i[7]^data_i[9]^data_i[10]^data_i[12]^data_i[13]^data_i[14]^data_i[15]^data_i[19]^data_i[21]^data_i[24]^data_i[26]^data_i[27]^data_i[34]^data_i[35]^data_i[39]^data_i[42]^data_i[43]^data_i[46]^data_i[50]^data_i[51]^data_i[53]^data_i[58]^data_i[59]^data_i[60];
  assign syndrome[7] = ecc_i[7]^data_i[1]^data_i[3]^data_i[4]^data_i[5]^data_i[6]^data_i[8]^data_i[9]^data_i[10]^data_i[13]^data_i[14]^data_i[15]^data_i[18]^data_i[20]^data_i[23]^data_i[25]^data_i[26]^data_i[31]^data_i[33]^data_i[34]^data_i[38]^data_i[41]^data_i[42]^data_i[45]^data_i[49]^data_i[50]^data_i[52]^data_i[57]^data_i[58]^data_i[59];

  //  clock has been gated in data_array
  always_ff @(posedge clk) begin
    syndrome_next <= syndrome;
    data_next     <= data_i;
  end

  always_comb begin
    error_mask = 64'b0;
    uncorrectable_error_o = 1'b0;
    unique case(syndrome_next)
      //  single error
      8'b00111011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001;
      8'b11101100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010;
      8'b01101110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100;
      8'b10011011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000;
      8'b11100110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000;
      8'b10111001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000;
      8'b11011100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000;
      8'b01000011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000;
      8'b10100111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000;
      8'b11101001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000;
      8'b11110100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000;
      8'b00111101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000;
      8'b01111100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000;
      8'b11110001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000;
      8'b11000111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000;
      8'b11111000: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000;
      8'b00111110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000;
      8'b00100101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000;
      8'b10010010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000;
      8'b01001001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000;
      8'b10100100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000;
      8'b01010010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000;
      8'b00101001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000;
      8'b10010100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000;
      8'b01001010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000;
      8'b10100001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000;
      8'b11010000: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000;
      8'b01101000: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000;
      8'b00110100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000;
      8'b00011010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000;
      8'b00001101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000;
      8'b10000110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000;
      8'b00100011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10010001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11001000: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01100100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00110010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00011001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10001100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01000110: error_mask = 64'b0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00010011: error_mask = 64'b0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10001001: error_mask = 64'b0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11000100: error_mask = 64'b0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01100010: error_mask = 64'b0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00110001: error_mask = 64'b0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10011000: error_mask = 64'b0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01001100: error_mask = 64'b0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00100110: error_mask = 64'b0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00001011: error_mask = 64'b0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10000101: error_mask = 64'b0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11000010: error_mask = 64'b0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01100001: error_mask = 64'b0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10110000: error_mask = 64'b0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01011000: error_mask = 64'b0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00101100: error_mask = 64'b0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00010110: error_mask = 64'b0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00000111: error_mask = 64'b0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10000011: error_mask = 64'b0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11000001: error_mask = 64'b0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11100000: error_mask = 64'b0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01110000: error_mask = 64'b0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00111000: error_mask = 64'b0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00011100: error_mask = 64'b0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00001110: error_mask = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      //  double adjacent error
      8'b11010111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011;
      8'b10000010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110;
      8'b11110101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100;
      8'b01111101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000;
      8'b01011111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000;
      8'b01100101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000;
      8'b10011111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000;
      8'b11100100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000;
      8'b01001110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000;
      8'b00011101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000;
      8'b11001001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000;
      8'b01000001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000;
      8'b10001101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000;
      8'b00110110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000;
      8'b00111111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000;
      8'b11000110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000;
      8'b00011011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000;
      8'b10110111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000;
      8'b11011011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000;
      8'b11101101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000;
      8'b11110110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000;
      8'b01111011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000;
      8'b10111101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000;
      8'b11011110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000;
      8'b11101011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000;
      8'b01110001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000;
      8'b10111000: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000;
      8'b01011100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000;
      8'b00101110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000;
      8'b00010111: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000;
      8'b10001011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000;
      8'b10100101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000;
      8'b10110010: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01011001: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10101100: error_mask = 64'b0000_0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01010110: error_mask = 64'b0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00101011: error_mask = 64'b0000_0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10010101: error_mask = 64'b0000_0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11001010: error_mask = 64'b0000_0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01010101: error_mask = 64'b0000_0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10011010: error_mask = 64'b0000_0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01001101: error_mask = 64'b0000_0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10100110: error_mask = 64'b0000_0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01010011: error_mask = 64'b0000_0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10101001: error_mask = 64'b0000_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11010100: error_mask = 64'b0000_0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01101010: error_mask = 64'b0000_0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00101101: error_mask = 64'b0000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10001110: error_mask = 64'b0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01000111: error_mask = 64'b0000_0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10100011: error_mask = 64'b0000_0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11010001: error_mask = 64'b0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b11101000: error_mask = 64'b0000_0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01110100: error_mask = 64'b0000_0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00111010: error_mask = 64'b0000_0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00010001: error_mask = 64'b0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10000100: error_mask = 64'b0000_0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01000010: error_mask = 64'b0000_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00100001: error_mask = 64'b0000_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b10010000: error_mask = 64'b0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b01001000: error_mask = 64'b0011_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00100100: error_mask = 64'b0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      8'b00010010: error_mask = 64'b1100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
      default: begin
        error_mask = 64'b0;
        uncorrectable_error_o = (syndrome == 64'b0) ? 1'b0 : 1'b1;
      end
    endcase
  end

  assign corrected_data_o = data_next ^ error_mask;

endmodule
